typedef enum {
		DIV,DIVU,REM,REMU
} ALU_func deriving(Eq, Bits, FShow);
