/*Copyright (c) 2013, IIT Madras
All rights reserved.

Redistribution and use in source and binary forms, with or without modification, are permitted provided that the following conditions are met:

*  Redistributions of source code must retain the above copyright notice, this list of conditions and the following disclaimer.
*  Redistributions in binary form must reproduce the above copyright notice, this list of conditions and the following disclaimer in the documentation and/or other materials provided with the distribution.
*  Neither the name of IIT Madras  nor the names of its contributors may be used to endorse or promote products derived from this software without specific prior written permission.

THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE. 
---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------

Module Name: RISCV 64bit Multiplier
Author Name: Rishi Naidu
Email id:    rishinaidu.rn@gmail.com
Last updated on : 11th October 2013

This is a pipelined integer multiplier that multiplies in five rg_clock cycles. 
Pipelining is implemented using FIFO registers in between the different stages of the multiplier.
This helps in improving the through put of the multiplier.

*********Performance****************:
Using UMCIP 65nm library in SYNOPSYS
Critical Path Length    :    0.5979 ns
Frequency 	        :    1.64 GHz
Combinational Cell Count:    57845
Sequential Cell Count   :    18810

Critical path : ff_stage1 ----> ff_stage2


******Refernce*******:
Redundant binary addition (IEEE paper "An 8.8-ns54 x 54-Bit Multiplier with High Speed Redundant Binary Architecture") 


The six stages of the multiplier are as follows

************Stage 1**************:

The Booth's 2nd algorithm is used to generate the partial products. Since the input size is 64 bits, the number of partial products generated is 32 (n/2). Alternate partial products are negated in order to generate redundant binary numbers. THis is unsigned booth multiplier, so an extra partial product is generated, which is due to zero extention of the multiplier.Two more partial products are used for Redundant binary addition. These partial products are then stored in the FIFO 'stage1'. Along with parameters to determine the type of multiplication instrcution.
************Stage 2***************:
Becoz of the high delay of RBA adder the addition of partial product take place in 3 stages.
The Redundant binary numbers are generated by grouping the i th and the (i+1)th partial products. Then these Redundant Binary Partial Products are added using a Wallace tree of redundant binary adders.
In stage2 16 partial products are added using RBA in 3 levels to generate a pair of RB number (RB_1)
The leaf of the wallace tree has 4 RB Adders that adds 8 RB numbers producing 4 RB numbers. These four RB numbers are the inputs to the 2 RB Adders in the next level of the wallace tree.The two RB number are in turn input to a final RBA adder to generate 1 pair of RB number. Next set of 16 partial products and extra partial product along with the result from stage 2 is stored in FIFO 'stage2'. Parameters to determine type of MUL instructions are also passed to next stage.

************Stage 3***************:
Input from FIFO 'stage2' includes the vector of partial products and the result of addition of 16 partial products.
In stage 3 next 16 partial products are added using RBA in 3 levels to generate a RB number(RB_2) (Same functions as in Stage2 is used)
RB_1 (generated in stage2) and RB_2 (generated in stage3) are stored in FIFO 'stage3', along with extra partial product and Parameters to determine type of MUL instructions are also passed to next stage.


************Stage 4***************:
The two rb number from FIFO 'stage3' are added along with a another rb number is added in 2 levels using RBA number.
level 1: RB_1 and RB_2
level 2: result from level 1 and another RB number (which is required to be added becoz of the logic in redundant binary adder)

The final RB number from stage 4 is stored in FIFO 'stage4' along with extra partial product and Parameters to determine type of MUL instructions are also passed to next stage.

************Stage 5***************:
The redundant binary product generated in the previous stage is converted into Normal Binary form by using RB to NB converter, then added to the extra partial product.The value is then passed to next stage using stage5 FIFO

************Stage6****************:
The value from FIFO stage5 is then converted to desired result based on the MUL type instruction. The resultant product is stored in the FIFO 'final_result'.

*/	




package integer_multiplier_riscv;

`include "defined_parameters.bsv"
import RB_NB::*;      //contain function to convert redundant binary number to normal binary number (Stage5)
import RBA::*;	      //contain functions for wallace tree redudant binary addition (Stage2,3,4)
import Booth2_pp_gen::*;//contain function to get partial products based on booth encoding (Stage1)
import Vector::*;
import FIFO::*;
import SpecialFIFOs::*;
import riscv_types::*;
//import decoder::*;

// The interface for the Integer Multiplier which accepts two 64 bit operands and produce 128 bit result
interface Ifc_integer_multiplier_riscv;

		/* Input Methods */
	method Action _start(Bit#(`REG_WIDTH) _in1, Bit#(`REG_WIDTH) _in2, ALU_func _mul_name,Bit#(1) _word_flag,  Bit#(TLog#(`TOTAL_THREADS)) thread_id, Bit#(TLog#(`PRF_SIZE)) _destination);// Start method to get inputs.
	method Action _set_flush(Bool _flush);   // Method to flush all FIFOs	
	method Action _release(); 		// Method to clear the result FIFO

		/* Output Methods */
	method Bit#(`REG_WIDTH) result_();	//Method to get result
	method Bit#(TLog#(`TOTAL_THREADS)) thread_id_();
	method Bit#(TLog#(`PRF_SIZE)) destination_address_();

endinterface:Ifc_integer_multiplier_riscv


/*
Following are the types of the structures used in each stage of the pipeline
*/
typedef struct{
	Vector#(TDiv#(`REG_WIDTH,2),Bit#(TMul#(`REG_WIDTH,2))) stage1; //Will store the 32 partial products generated in stage1
	Bit#(2) stage1_mul_type;     // TO determine the type of MUL instruction to be used in last stage to get final 64  bit result
	Bit#(1) stage1_word_flag;    // To determine if its a word instruction or not to be used in last stage to get final 64 bit result
	Bit#(1) stage1_sign_bit_op1; // Operand1 sign bit to be used in last stage to get final 64 bit result                            
	Bit#(1) stage1_sign_bit_op2; // Operand2 sign bit to be used in last stage to get final 64 bit result  
	Bit#(TMul#(`REG_WIDTH,2)) stage1_extra_pp;   //Generated due to Unsigned multiplication in booth                   
	Bit#(TLog#(`TOTAL_THREADS)) thread_id;
	Bit#(TLog#(`PRF_SIZE)) destination;	// destination address where the output is to be written in the Regfile
}Stage1_data deriving(Eq,Bits);

typedef struct{
	Bit#(TMul#(`REG_WIDTH,4)) data_computed_stage2; //Will store result of addition of 16 partial products computed in stage2
	Vector#(TDiv#(`REG_WIDTH,4),Bit#(TMul#(`REG_WIDTH,2))) vector_pp; // Will again store the 32 partial products passed from stage1
	Bit#(2) stage2_mul_type;        // TO determine the type of MUL instruction to be used in last stage to get final 64  bit result
	Bit#(1) stage2_word_flag;       // To determine if its a word instruction or not to be used in last stage to get final 64 bit result
	Bit#(1) stage2_sign_bit_op1;    // Operand1 sign bit to be used in last stage to get final 64 bit result                            
	Bit#(1) stage2_sign_bit_op2;    // Operand2 sign bit to be used in last stage to get final 64 bit result                            
	Bit#(TMul#(`REG_WIDTH,2)) stage2_extra_pp;      //Generated due to Unsigned multiplication in booth                   
	Bit#(TLog#(`TOTAL_THREADS)) thread_id;
	Bit#(TLog#(`PRF_SIZE)) destination;	// destination address where the output is to be written in the Regfile
}Stage2_data deriving(Eq,Bits);

typedef struct{
	Bit#(TMul#(`REG_WIDTH,4)) data_from_stage2; //Will store result of addition of 1st set of 16 partial products
	Bit#(TMul#(`REG_WIDTH,4)) data_from_stage3; //Will store result of addition of 2nd set of 16 partial products
	Bit#(2) stage3_mul_type;        // TO determine the type of MUL instruction to be used in last stage to get final 64  bit result
	Bit#(1) stage3_word_flag;       // To determine if its a word instruction or not to be used in last stage to get final 64 bit result
	Bit#(1) stage3_sign_bit_op1;    // Operand1 sign bit to be used in last stage to get final 64 bit result                            
	Bit#(1) stage3_sign_bit_op2;    // Operand2 sign bit to be used in last stage to get final 64 bit result                            
	Bit#(TMul#(`REG_WIDTH,2)) stage3_extra_pp;       //Generated due to Unsigned multiplication in booth                   
	Bit#(TLog#(`TOTAL_THREADS)) thread_id;
	Bit#(TLog#(`PRF_SIZE)) destination;	// destination address where the output is to be written in the Regfile
}Stage3_data deriving(Eq,Bits);

typedef struct{
	Bit#(TMul#(`REG_WIDTH,4)) final_rb_number; //Will store the final RB number computed in stage4
	Bit#(2) stage4_mul_type;      // TO determine the type of MUL instruction to be used in last stage to get final 64  bit result
	Bit#(1) stage4_word_flag;     // To determine if its a word instruction or not to be used in last stage to get final 64 bit result
	Bit#(1) stage4_sign_bit_op1;  // Operand1 sign bit to be used in last stage to get final 64 bit result                            
	Bit#(1) stage4_sign_bit_op2;  // Operand2 sign bit to be used in last stage to get final 64 bit result                            
	Bit#(TMul#(`REG_WIDTH,2)) stage4_extra_pp;        //Generated due to Unsigned multiplication in booth                   
	Bit#(TLog#(`TOTAL_THREADS)) thread_id;
	Bit#(TLog#(`PRF_SIZE)) destination;	// destination address where the output is to be written in the Regfile

}Stage4_data deriving(Eq,Bits);


typedef struct{ 
	Bit#(TMul#(`REG_WIDTH,2)) unsigned_mul_output; // Unsigned multiplication after Rb to Nb conversion
	Bit#(2) stage5_mul_type;      // TO determine the type of MUL instruction to be used in last stage to get final 64  bit result
	Bit#(1) stage5_word_flag;     // To determine if its a word instruction or not to be used in last stage to get final 64 bit result
	Bit#(1) stage5_sign_bit_op1;  // Operand1 sign bit to be used in last stage to get final 64 bit result                            
	Bit#(1) stage5_sign_bit_op2;  // Operand2 sign bit to be used in last stage to get final 64 bit result                            
	Bit#(TLog#(`TOTAL_THREADS)) thread_id;
	Bit#(TLog#(`PRF_SIZE)) destination;	// destination address where the output is to be written in the Regfile
}Stage5_data deriving(Eq,Bits);


(*synthesize*)
module mkinteger_multiplier_riscv(Ifc_integer_multiplier_riscv);
	
	Wire#(Bool) wr_flush <-mkDWire(False);	 //Wire for flush
	FIFO#(Stage1_data) ff_stage1 <- mkFIFO;  //This FIFO stores the 32 128 bit partial products produced in stage 1
	FIFO#(Stage2_data) ff_stage2 <- mkFIFO;	 //This FIFO stores the result of addition of 1st set of 16 partial products and the 32 128 bit partial products computed in stage1
	FIFO#(Stage3_data) ff_stage3 <- mkFIFO;	 //This FIFO stores the result of the 1st set and 2nd set of 16 partial products computed in stage 2 and 3 respectively
	FIFO#(Stage4_data) ff_stage4 <- mkFIFO;	 //This FIFO stores the result of the Redundant Binary Addition of the Redundant Binary Partial Products
	FIFO#(Stage5_data) ff_stage5 <- mkFIFO;	 //This FIFO stores the normal binary product after conversion from rb number	
	FIFO#(Bit#(`REG_WIDTH)) ff_final_result <- mkBypassFIFO;	 //This FIFO stores the final 64 bit result of MUL instructions
	Reg#(Bool) rg_ready_signal <-mkReg(False);
	Reg#(Bit#(TLog#(`TOTAL_THREADS))) rg_thread_id <-mkReg(0);
	FIFO#(Bit#(TLog#(`PRF_SIZE))) ff_destination_address<-mkBypassFIFO();
	/* This rule is fired only when the wr_flush signal is invoked.
	Here all the fifos are cleared and thus any comutation is abandoned.
	*/
	rule rl_flush_data(wr_flush);
		ff_stage1.clear();
		ff_stage2.clear();
		ff_stage3.clear();
		ff_stage4.clear();
	    ff_stage5.clear();
		ff_final_result.clear();
		ff_destination_address.clear();
		rg_ready_signal<=False; // False when flusshed
		rg_thread_id<=0;
	endrule:rl_flush_data
	

	//Stage 2
	rule rl_wallace_tree_part1(!wr_flush);
		//$display("Executing Integer MUL stage 2"); 
		let lv_data_stage1=ff_stage1.first;    //Get the 32 partial products from FIFO stage1
		ff_stage1.deq;	
		Vector#(TDiv#(`REG_WIDTH,4),Bit#(TMul#(`REG_WIDTH,2))) upper_half = take(lv_data_stage1.stage1);
		let lv_result_stage2=wallace_rba(upper_half);
		
		ff_stage2.enq(Stage2_data{data_computed_stage2:lv_result_stage2, //Forward result to next stage
					vector_pp:takeTail(lv_data_stage1.stage1), //Forward the 32 partial product for addition of next 16 partial products in stage3
					stage2_mul_type:     lv_data_stage1.stage1_mul_type,
					stage2_word_flag:    lv_data_stage1.stage1_word_flag,
					stage2_sign_bit_op1: lv_data_stage1.stage1_sign_bit_op1,
					stage2_extra_pp: lv_data_stage1.stage1_extra_pp,
					thread_id:lv_data_stage1.thread_id,
					destination:lv_data_stage1.destination,
					stage2_sign_bit_op2: lv_data_stage1.stage1_sign_bit_op2});

	endrule:rl_wallace_tree_part1

	//Stage 3
	rule rl_wallace_tree_part2(!wr_flush);
		//$display("Executing Integer MUL stage 3");
		let lv_data_stage2=ff_stage2.first;	//Get result of additon of 16 pp and the 32 pp's for next step of addition
//		Vector#(TDiv#(`REG_WIDTH,4),Bit#(TMul#(`REG_WIDTH,2))) lower_half = takeTail(lv_data_stage2.vector_pp);
		let lv_result_stage3= wallace_rba(lv_data_stage2.vector_pp);
		ff_stage2.deq;

		ff_stage3.enq(Stage3_data{data_from_stage2: lv_data_stage2.data_computed_stage2, //Result of additon of 1st 16 partial products
					  data_from_stage3: lv_result_stage3,      //Result of addition of next 16 partial products
					  stage3_mul_type:     lv_data_stage2.stage2_mul_type,
					  stage3_word_flag:    lv_data_stage2.stage2_word_flag,
					  stage3_sign_bit_op1: lv_data_stage2.stage2_sign_bit_op1,
					  stage3_extra_pp: lv_data_stage2.stage2_extra_pp,
					  thread_id:lv_data_stage2.thread_id, 
					destination:lv_data_stage2.destination,
					  stage3_sign_bit_op2: lv_data_stage2.stage2_sign_bit_op2
					});
	endrule:rl_wallace_tree_part2
	//Stage 4
	rule rl_wallace_tree_final(!wr_flush);
		//$display("Executing Integer MUL stage 4");
		let lv_data_stage3=ff_stage3.first;		// Get result of additon of both 1st 16 pp and next 16 pp
		let lv_result_stage4=wallace_rba_final(lv_data_stage3.data_from_stage2,lv_data_stage3.data_from_stage3); // Final RB number. An extra RB number is added in function due to logic in redundant binary addition
		ff_stage3.deq;

		ff_stage4.enq(Stage4_data{final_rb_number:lv_result_stage4,
					stage4_extra_pp: lv_data_stage3.stage3_extra_pp,		
					  stage4_mul_type:     lv_data_stage3.stage3_mul_type,
					  stage4_word_flag:    lv_data_stage3.stage3_word_flag,
					  stage4_sign_bit_op1: lv_data_stage3.stage3_sign_bit_op1,
					  thread_id:lv_data_stage3.thread_id,
					destination:lv_data_stage3.destination,
					  stage4_sign_bit_op2: lv_data_stage3.stage3_sign_bit_op2});  //FInal RB number in Stage 4 FIFO
	endrule:rl_wallace_tree_final



	//Stage5

	rule rl_rb_nb(!wr_flush);
		// The Redundant Binary product generated in the previous stage is converted into the normal binary form.
		
		let lv_data_stage4= ff_stage4.first(); // Get RB number generated in stage 4
//		let normal_binary_product=rb_nb(lv_data_stage4.final_rb_number) + lv_data_stage4.stage4_extra_pp; // Converted RB number is added to extra pp to get the final result of unsigned multiplication
//		let normal_binary_product = lv_data_stage4.final_rb_number[255:128] + (~lv_data_stage4.final_rb_number[127:0] +1)+lv_data_stage4.stage4_extra_pp;
		let normal_binary_product = lv_data_stage4.final_rb_number[(`REG_WIDTH*4)-1:(`REG_WIDTH*2)] + (~lv_data_stage4.final_rb_number[(`REG_WIDTH*2)-1:0] +1)+lv_data_stage4.stage4_extra_pp;
		ff_stage4.deq();
		
		ff_stage5.enq(Stage5_data{unsigned_mul_output : normal_binary_product,		
					  stage5_mul_type:     lv_data_stage4.stage4_mul_type,
					  stage5_word_flag:    lv_data_stage4.stage4_word_flag,
					  stage5_sign_bit_op1: lv_data_stage4.stage4_sign_bit_op1,
					  thread_id:lv_data_stage4.thread_id,
					destination:lv_data_stage4.destination,
					  stage5_sign_bit_op2: lv_data_stage4.stage4_sign_bit_op2 });
	
	endrule:rl_rb_nb
	
	//Stage6
	rule rl_final_output(!wr_flush);
		//Changing the final answer based on different multiplier instruction, before storing in final_result FIFO
		// _mul_type  determines if its MUL, MULH, MULHSU, MULHU
		//_word_flag determines if its MULW instruction or not
		let lv_data_stage5 = ff_stage5.first();
		rg_thread_id<=lv_data_stage5.thread_id;
		ff_destination_address.enq(lv_data_stage5.destination);
		Bit#(TMul#(`REG_WIDTH,2)) unsigned_output = lv_data_stage5.unsigned_mul_output; 
		ff_stage5.deq;
		Bit#(`REG_WIDTH) _final_result= 0;

		`ifdef Multiplier64	
			if (lv_data_stage5.stage5_word_flag==1) begin //MULW
				_final_result = signExtend(unsigned_output[31:0]);	
			end
			else begin

				case (lv_data_stage5.stage5_mul_type) matches
					2'b00: begin//MUL (Simple MUL,output is lower 64 bits)
						_final_result = unsigned_output[`REG_WIDTH-1:0];
					end
					2'b01: begin//MULH (SignedxSigned Multiplication output is higher 64 bits)
						Bit#(TMul#(`REG_WIDTH,2)) lv_result_temp = ((lv_data_stage5.stage5_sign_bit_op1^lv_data_stage5.stage5_sign_bit_op2)==1) ? (~unsigned_output + 1): unsigned_output ;	
						_final_result = lv_result_temp[(`REG_WIDTH*2)-1:`REG_WIDTH];
					end
					2'b10: begin//MULHSU (SignedxUnsigned Multiplication output is higher 64 bits)
						Bit#(TMul#(`REG_WIDTH,2)) lv_temp_result = (lv_data_stage5.stage5_sign_bit_op1==1) ? (~unsigned_output + 1): unsigned_output ;
						_final_result = lv_temp_result[(`REG_WIDTH*2)-1:`REG_WIDTH];
					end
					2'b11: begin//MULHU (Unsigned Multiplication, output is higher 64 bits)
						_final_result = unsigned_output[(`REG_WIDTH*2)-1:`REG_WIDTH];
					end

				endcase
			end
		`else
				case (lv_data_stage5.stage5_mul_type) matches
					2'b00: begin//MUL (Simple MUL,output is lower 64 bits)
						_final_result = unsigned_output[`REG_WIDTH-1:0];
					end
					2'b01: begin//MULH (SignedxSigned Multiplication output is higher 64 bits)
						Bit#(TMul#(`REG_WIDTH,2)) lv_result_temp = ((lv_data_stage5.stage5_sign_bit_op1^lv_data_stage5.stage5_sign_bit_op2)==1) ? (~unsigned_output + 1): unsigned_output ;	
						_final_result = lv_result_temp[(`REG_WIDTH*2)-1:`REG_WIDTH];
					end
					2'b10: begin//MULHSU (SignedxUnsigned Multiplication output is higher 64 bits)
						Bit#(TMul#(`REG_WIDTH,2)) lv_temp_result = (lv_data_stage5.stage5_sign_bit_op1==1) ? (~unsigned_output + 1): unsigned_output ;
						_final_result = lv_temp_result[(`REG_WIDTH*2)-1:`REG_WIDTH];
					end
					2'b11: begin//MULHU (Unsigned Multiplication, output is higher 64 bits)
						_final_result = unsigned_output[(`REG_WIDTH*2)-1:`REG_WIDTH];
					end

				endcase
		`endif


		ff_final_result.enq(_final_result);  //  Normal binary product stored in the final result FIFO
		//$display("Executing Integer MUL stage 5. Output=%h",_final_result); 
	
		rg_ready_signal <=True; // Assign ready Signal TRUE, as result is available
	endrule:rl_final_output

	method Action _start(Bit#(`REG_WIDTH) _in1, Bit#(`REG_WIDTH) _in2, ALU_func _mul_name,Bit#(1) _word_flag,  Bit#(TLog#(`TOTAL_THREADS)) thread_id, Bit#(TLog#(`PRF_SIZE)) _destination) if(!wr_flush);
		Bit#(`REG_WIDTH) _operand1 = 0;
		Bit#(`REG_WIDTH) _operand2 = 0;
		Bit#(1) _sign_bit_op2 = _in2[`REG_WIDTH-1];  // Sign bit operand1 for propogation across different stages to be used in the final stage
		Bit#(1) _sign_bit_op1 = _in1[`REG_WIDTH-1];  //Sign bit operand1 for propogation across different stages to be used in the final stage
		Bit#(2) _mul_type = 0;

		case (_mul_name)
			MUL : 	_mul_type = 'b00;
			MULH: 	_mul_type = 'b01;
			MULHSU:	_mul_type = 'b10;
			MULHU:  _mul_type = 'b11;
			//MULW : 	_mul_type = 'b100;
			//MULHW: 	_mul_type = 'b101;
			//MULHSUW:_mul_type = 'b110;
			//MULHUW: _mul_type = 'b111;			
		endcase
				
		// Changing operand1 and operand2 based on different multiplier instruction before feeding it into the multiplier module
		// _mul_type  determines if its MUL, MULH, MULHSU, MULHU
		//_word_flag determines if its MULW instruction or not
		`ifdef Multiplier64
			if (_word_flag==1) begin //MULW (Word instruction, multiplication of lower 32 bits where output is signextended lower 32 bits output)
				_operand1 = {32'b0,_in1[31:0]};
				_operand2 = {32'b0,_in2[31:0]};
			end
			else begin

				if((_mul_type[0]^_mul_type[1])==0)
					_operand1 = _in1;
				else
					_operand1 = _in1[`REG_WIDTH-1]==1? (~_in1 +1) :_in1;

				if(_mul_type==2'b01)
					_operand2=_in2[`REG_WIDTH-1]==1? (~_in2 +1) :_in2;
				else
					_operand2=_in2;

			end
		`else
				if((_mul_type[0]^_mul_type[1])==0)
					_operand1 = _in1;
				else
					_operand1 = _in1[`REG_WIDTH-1]==1? (~_in1 +1) :_in1;

				if(_mul_type==2'b01)
					_operand2=_in2[`REG_WIDTH-1]==1? (~_in2 +1) :_in2;
				else
					_operand2=_in2;
		`endif
		$display("_operand1 = %h , _operand2 = %h", _operand1,_operand2);
		Bit#(TAdd#(`REG_WIDTH,3)) lv_mult={2'b00,_operand1,0};		// lv_mult     = multiplier appended with a zero and extended with zeros, a requirement of booth's unsigned multiplication of second order algorithm
		Bit#(TMul#(`REG_WIDTH,2)) lv_multp=zeroExtend(_operand2);	// lv_multp    = multiplicand
                
	
		Bit#(TMul#(`REG_WIDTH,2)) lv_lmultp = lv_multp<<1;	// lv_lmultp    = multiplicand left shifted one bit position/ twice of multiplicand requied for booth encoding
			
		// Generation of the 32 partial products using Booth's second order algorithm. The i+1 i i-1 th bits are used as the select bits
		// These 32 partial products are converted into redundant binary partial products by taking two at a time.i.e every adjacent partial product.
		// To form a RB number, the two's complement of the second number is needed. So, every odd numbered partial product is inverted. To avoid an addition of 1
		// which will involve a a carry propagation, we take these 16 1's along with a 128'b0 to form the 9th partial product.
		// The last two bit positions is due to the left shifting of two bits for adjacent partial products. Since, the odd numbered partial products
		// are inverted, we append one's. For even numbered partial products, we append zeroes.
		
		Vector#(TDiv#(`REG_WIDTH,2),Bit#(TMul#(`REG_WIDTH,2))) lv_pp = replicate(0); // Creating a vector for 32 128 bit pp's
		Bit#(TMul#(`REG_WIDTH,2)) lv_extra_pp = 0; //Extra partial product generated due to the 2 zero bit extended in multiplier for unsigned multiplication
		lv_pp[0]=gen_pp (lv_multp,lv_lmultp,lv_mult[2:0],0);
		lv_pp[1]=(gen_pp(lv_multp,lv_lmultp,lv_mult[4:2],1)<<2 | 'b11);
		lv_pp[2]=(gen_pp(lv_multp,lv_lmultp,lv_mult[6:4],0)<<4);
		lv_pp[3]=(gen_pp(lv_multp,lv_lmultp,lv_mult[8:6],1)<<2 | 'b11)<<4;
		
		`ifdef Multiplier16
			lv_pp[4]=(gen_pp(lv_multp,lv_lmultp,lv_mult[10:8],0)<<8);
			lv_pp[5]=(gen_pp(lv_multp,lv_lmultp,lv_mult[12:10],1)<<2 | 'b11)<<8;
			lv_pp[6]=(gen_pp(lv_multp,lv_lmultp,lv_mult[14:12],0)<<12);
			lv_pp[7]=(gen_pp(lv_multp,lv_lmultp,lv_mult[16:14],1)<<2 | 'b11)<<12;
		`endif

		`ifdef Multiplier32
			lv_pp[8]=(gen_pp(lv_multp,lv_lmultp,lv_mult[18:16],0)<<16);
			lv_pp[9]=(gen_pp(lv_multp,lv_lmultp,lv_mult[20:18],1)<<2 | 'b11)<<16;
			lv_pp[10]=(gen_pp(lv_multp,lv_lmultp,lv_mult[22:20],0)<<20);
			lv_pp[11]=(gen_pp(lv_multp,lv_lmultp,lv_mult[24:22],1)<<2 | 'b11)<<20;
			lv_pp[12]=(gen_pp(lv_multp,lv_lmultp,lv_mult[26:24],0)<<24);
			lv_pp[13]=(gen_pp(lv_multp,lv_lmultp,lv_mult[28:26],1)<<2 | 'b11)<<24;
			lv_pp[14]=(gen_pp(lv_multp,lv_lmultp,lv_mult[30:28],0)<<28);
			lv_pp[15]=(gen_pp(lv_multp,lv_lmultp,lv_mult[32:30],1)<<2 | 'b11)<<28;
		`endif
 
		`ifdef Multiplier64
			lv_pp[16]=(gen_pp(lv_multp,lv_lmultp,lv_mult[34:32],0)<<32);
			lv_pp[17]=(gen_pp(lv_multp,lv_lmultp,lv_mult[36:34],1)<<2 | 'b11)<<32;
			lv_pp[18]=(gen_pp(lv_multp,lv_lmultp,lv_mult[38:36],0)<<36);
			lv_pp[19]=(gen_pp(lv_multp,lv_lmultp,lv_mult[40:38],1)<<2 | 'b11)<<36;
			lv_pp[20]=(gen_pp(lv_multp,lv_lmultp,lv_mult[42:40],0)<<40);
			lv_pp[21]=(gen_pp(lv_multp,lv_lmultp,lv_mult[44:42],1)<<2 | 'b11)<<40;
			lv_pp[22]=(gen_pp(lv_multp,lv_lmultp,lv_mult[46:44],0)<<44);
			lv_pp[23]=(gen_pp(lv_multp,lv_lmultp,lv_mult[48:46],1)<<2 | 'b11)<<44;
			lv_pp[24]=(gen_pp(lv_multp,lv_lmultp,lv_mult[50:48],0)<<48);
			lv_pp[25]=(gen_pp(lv_multp,lv_lmultp,lv_mult[52:50],1)<<2 | 'b11)<<48;
			lv_pp[26]=(gen_pp(lv_multp,lv_lmultp,lv_mult[54:52],0)<<52);
			lv_pp[27]=(gen_pp(lv_multp,lv_lmultp,lv_mult[56:54],1)<<2 | 'b11)<<52;
			lv_pp[28]=(gen_pp(lv_multp,lv_lmultp,lv_mult[58:56],0)<<56);
			lv_pp[29]=(gen_pp(lv_multp,lv_lmultp,lv_mult[60:58],1)<<2 | 'b11)<<56;
			lv_pp[30]=(gen_pp(lv_multp,lv_lmultp,lv_mult[62:60],0)<<60);
			lv_pp[31]=(gen_pp(lv_multp,lv_lmultp,lv_mult[64:62],1)<<2 | 'b11)<<60;
			lv_extra_pp[127:64] = gen_pp(lv_multp,lv_lmultp,lv_mult[66:64],0)[63:0];
		`endif

		
		// The 32 partial products are stored in the stage1 FIFO along with parameters to determine MUL type and the extra pp
		ff_stage1.enq(Stage1_data{stage1:lv_pp,// Storing the partial products in the final FIFO
					stage1_extra_pp : lv_extra_pp,
					stage1_mul_type: _mul_type,stage1_word_flag: _word_flag, 
					thread_id:thread_id,
					destination: _destination,
					stage1_sign_bit_op1: _sign_bit_op1,stage1_sign_bit_op2:_sign_bit_op2}); 
	endmethod


	method Bit#(`REG_WIDTH) result_();   //Method to get the result
		return ff_final_result.first;
	endmethod
	
	method Action _set_flush(Bool _flush); // Method to flush the pipe
		wr_flush<=_flush;
	endmethod

	method Action _release(); // Method to release the final result FIFO after obtaining result
		ff_final_result.deq();
		ff_destination_address.deq();
	endmethod

	
	method Bit#(TLog#(`TOTAL_THREADS)) thread_id_();
		return rg_thread_id;
	endmethod
	method Bit#(TLog#(`PRF_SIZE)) destination_address_();
		return ff_destination_address.first();
	endmethod
endmodule:mkinteger_multiplier_riscv

endpackage:integer_multiplier_riscv
