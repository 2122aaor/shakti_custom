/*


-------------------------------------------------------------------------------
-- 
-- Copyright (C) 2013 Indian Institute of Technology Madras (IITM)
-- All rights reserved.
-- 
-- This source file may be used and distributed without
-- restriction provided that this copyright statement is not
-- removed from the file and that any derivative work contains
-- the original copyright notice and the associated disclaimer.
-- 
-- This source file is free software; you can redistribute it
-- and/or modify it under the terms of the GNU General
-- Public License as published by the Free Software Foundation;
-- either version 3.0 of the License, or (at your option) any
-- later version.
-- 
-- 
-- You should have received a copy of the GNU General
-- Public License along with this source;
--
-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDER ``AS IS'' AND ANY EXPRESS
-- OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES
-- OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN
-- NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE FOR ANY
-- DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
-- LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND
-- ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
-- (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF
-- THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
--
-- The views and conclusions contained in the software and documentation are
-- those of the authors and should not be interpreted as representing official
-- policies, either expressed or implied, of the copyright holder.
-- 
-------------------------------------------------------------------------------


Module Name: Interger Multiplier used in Floating Point Unit.
Author Name: Neel Gala , Kalyan Kumar, Aditya Govardhan, Vinod.G
Email Id: neelgala@gmail.com kalyavkumar.suvvada@gmail.com, dtgovardhan@gmail.com, g.vinod1993@gmail.com
Last updated on : 30th September, 2013

This is a pipelined integer multiplier that multiplies in four clock cycles. 
Pipelining is implemented using FIFO registers in between the different stages of the multiplier.
This helps in improving the through put of the multiplier.

The Four stages of the multiplier are as follows

Stage 1:

The Booth's 2nd algorithm is used to generate the partial products. Since the input size is 32 bits, the number of partial products generated is 16. Alternate partial products are negated in order to generate redundant binary numbers. Two more partial products are used for Redundant binary addition. These partial products are then stored in the FIFO 'stage2'.

Stage 2:

The Redundant binary numbers are generated by grouping the i th and the (i+1)th partial products. Then these Redundant Binary Partial Products are added using a Wallace tree of redundant binary adders.Due to the high delay of the RB Adders, the wallace tree multiplication is split into two cycles.

The leaf of the wallace tree has 4 RB Adders that adds 8 RB numbers producing 4 RB numbers. These four RB numbers are the inputs to the 2 RB Adders in the next level of the wallace tree. Finally, this stage produces 2 RB. Now, totally we have added 8 RB numbers. We still have 1 un_added RB number and two results produced from this stage.

Stage 3
 These 3 RB numbers are added with a 2 level RB Adder with one RB Adder in each level. This stage finally produces the result of the addition process. The result, also a redundant binary number, is stored in the FIFO 'stage3'.

Stage 4

The redundant binary product generated in the previous stage is converted into Normal Binary form by using RB to NB converter. The resultant product is stored in the FIFO 'prod'.

*/

package integermultiplier_for_spfpu;

import RB_NB::*;
import RBA::*;
import Vector::*;
import FIFO::*;


// Function to generate the Booth's partial products.
(*noinline*)
function Bit#(64) gen_pp(Bit#(64) multp, Bit#(64) lmultp, Bit#(3) sel, int inv);
	
	Bit#(64) result='d0;
	case(sel)
		'd0: result=64'b0; 	//zero
		'd1: result=multp; 	// M
		'd2: result=multp; 	// M
		'd3: result=lmultp;	// 2M
		'd4: result=~lmultp+1;	// -2M			
		'd5: result=~multp+1;	// -M
		'd6: result=~multp+1;	// -M
		'd7: result=64'b0;	// zero
	endcase

	//This inversion of alternate partial products is to obtain the redundant binary numbers from this and the previous partial product.
	if(inv==1)
		result=~result;
	
	return result;

endfunction


// The interface for the Integer Multiplier which accepts 2 32 bit operands(signed) and produces the 64 bit product as the output
interface Ifc_integer_multiplier_for_spfmul;
		/* Input Methods */
	method Action _start( Bit#(32) _operand1, Bit#(32) _operand2 , Bit#(32) _fsr, Bit#(3) rounding_mode, bit _sign, Bit#(10) _summed_exponent, bit _invalid, Bit#(1) _infinity, Bit#(1) _zero);
	method Action _deque();

		/* Output Methods */
	method Stage4_data result_();
endinterface:Ifc_integer_multiplier_for_spfmul

typedef struct{
	Bit#(32) fsr;			// the input fsr
    Bit#(3) rounding_mode;          // static rounding mode encoded in the instruction
	Bit#(10) summed_exponent;	// the sum of the exponents
	bit sign;			// the sign bit
	Bit#(1) infinity;		// the infinity Flag
	Bit#(1) invalid;		// the Invalid Flag
	Bit#(1) zero;			// The Zero Flag
	Vector#(16,Bit#(64)) stage1;	// partial product array.
	}Stage1_data deriving(Eq,Bits);

typedef struct{
	Bit#(32) fsr;                   // the input fsr
    Bit#(3) rounding_mode;          // static rounding mode encoded in the instruction
	Bit#(10) summed_exponent;	// the sum of the exponents.
	bit sign;			// the sign bit of the result
	Bit#(1) infinity;		// the infinity Flag
	Bit#(1) invalid;                // the Invalid Flag
	Bit#(1) zero;                   // The Zero Flag
	Bit#(384) stage2;
	}Stage2_data deriving(Eq,Bits);

typedef struct{
	Bit#(32) fsr;                   // the input fsr
    Bit#(3) rounding_mode;          // static rounding mode encoded in the instruction
	Bit#(10) summed_exponent;	// the sum of the exponents.
	bit sign;			// the sign bit of the result
	Bit#(1) infinity;		// the infinity Flag
	Bit#(1) invalid;                // the Invalid Flag
	Bit#(1) zero;                   // The Zero Flag
	Bit#(128) stage3;
	}Stage3_data deriving(Eq,Bits);

typedef struct{
	Bit#(32) fsr;                   // the input fsr
    Bit#(3) rounding_mode;          // static rounding mode encoded in the instruction
	Bit#(10) summed_exponent;	// the sum of the exponents.
	bit sign;			// the sign bit of the result
	Bit#(1) infinity;		// the infinity Flag
	Bit#(1) invalid;                // the Invalid Flag
	Bit#(1) zero;                   // The Zero Flag
	Bit#(145) stage3a;
	}Stage3a_data deriving(Eq,Bits);

typedef struct{
	Bit#(32) fsr;                   // the input fsr
    Bit#(3) rounding_mode;          // static rounding mode encoded in the instruction
	Bit#(10) summed_exponent;	// the sum of the exponents.
	bit sign;			// the sign bit of the result
	Bit#(1) infinity;		// the infinity Flag
	Bit#(1) invalid;                // the Invalid Flag
	Bit#(1) zero;                   // The Zero Flag
	Bit#(161) stage3b;
	}Stage3b_data deriving(Eq,Bits);

typedef struct{
	Bit#(32) fsr;                   // the input fsr
    Bit#(3) rounding_mode;          // static rounding mode encoded in the instruction
	Bit#(10) summed_exponent;	// the sum of the exponents.
	bit sign;			// the sign bit of the result
	Bit#(1) infinity;		// the infinity Flag
	Bit#(1) invalid;                // the Invalid Flag
	Bit#(1) zero;                   // The Zero Flag
	Bit#(177) stage3c;
	}Stage3c_data deriving(Eq,Bits);

typedef struct{
	Bit#(32) fsr;                   // the input fsr
    Bit#(3) rounding_mode;          // static rounding mode encoded in the instruction
	Bit#(10) summed_exponent;	// the sum of the exponents.
	bit sign;			// the sign bit of the result
	Bit#(1) infinity;		// the infinity Flag
	Bit#(1) invalid;                // the Invalid Flag
	Bit#(1) zero;                   // The Zero Flag
	Bit#(64) final_result;
	}Stage4_data deriving(Eq,Bits);



(*synthesize*)
module mkinteger_multiplier_for_spfmul(Ifc_integer_multiplier_for_spfmul);

	FIFO#(Stage1_data) ff_stage1 <- mkFIFO;  //This FIFO stores the 16 64 bit partial products produced in the previous cycle
	FIFO#(Stage2_data) ff_stage2 <- mkFIFO;	 //This FIFO stores the 3 Redundant binary numbers left to be added.3x2x64=384 bits
	FIFO#(Stage3_data) ff_stage3 <- mkFIFO;	 //This FIFO stores the result of the Redundant Binary Addition of the Redundant Binary Partial Products
	FIFO#(Stage3a_data) ff_stage3a <- mkFIFO;	 //This FIFO stores the result of the Redundant Binary Addition of the Redundant Binary Partial Products
	FIFO#(Stage3b_data) ff_stage3b <- mkFIFO;	 //This FIFO stores the result of the Redundant Binary Addition of the Redundant Binary Partial Products
	FIFO#(Stage3c_data) ff_stage3c <- mkFIFO;	 //This FIFO stores the result of the Redundant Binary Addition of the Redundant Binary Partial Products
	FIFO#(Stage4_data) ff_final_result <- mkFIFO;//This FIFO stores the result of the multiplication of the two operands after converting the RB number to NB

	//Cycle 2
	rule rl_wallace_tree_part1;
		//$display("Executing FMUL stage 2-1");
		// The first two levels of wallace tree addition is performed
		let lv_info1=ff_stage1.first;
		ff_stage1.deq;
		let lv_res=wallace_rba_part1(lv_info1.stage1);
		let lv_s2_1p=lv_res[255:192];
		let lv_s2_1m=lv_res[191:128];
		let lv_s2_2p=lv_res[127:64];
		let lv_s2_2m=lv_res[63:0];
		// The 3 redundant binary partial products, 2 from the result of this stage and one from the previous stage.
		ff_stage2.enq(Stage2_data{
									fsr:lv_info1.fsr,
				                    rounding_mode : lv_info1.rounding_mode,
									summed_exponent:lv_info1.summed_exponent,
									sign : lv_info1.sign,
									infinity:lv_info1.infinity,
									invalid:lv_info1.invalid,
									zero:lv_info1.zero,
									stage2:{lv_info1.stage1[14],lv_info1.stage1[15],lv_s2_1p,lv_s2_1m,lv_s2_2p,lv_s2_2m}
					});
	endrule:rl_wallace_tree_part1

	//cycle 3
	rule rl_wallace_tree_part2;
		//$display("Executing FMUL stage 2-2");
		// The addition of the remaining 3 RB Numbers is completed in this stage.
		let lv_info2=ff_stage2.first;
		let lv_inp1=lv_info2.stage2[383:320];
		let lv_inp2=lv_info2.stage2[319:256];
		let lv_s2_1p=lv_info2.stage2[255:192];
		let lv_s2_1m=lv_info2.stage2[191:128];
		let lv_s2_2p=lv_info2.stage2[127:64];
		let lv_s2_2m=lv_info2.stage2[63:0];
		ff_stage2.deq;
		// Res is the required product of the two operands but in the redundant binary format
		let lv_res=wallace_rba_part2(lv_s2_1p,lv_s2_1m,lv_s2_2p,lv_s2_2m,lv_inp1,lv_inp2);
		ff_stage3.enq(Stage3_data{
									fsr:lv_info2.fsr,
				                    rounding_mode : lv_info2.rounding_mode,
									summed_exponent:lv_info2.summed_exponent,
									sign : lv_info2.sign,
									infinity:lv_info2.infinity,
									invalid:lv_info2.invalid,
									zero:lv_info2.zero,
									stage3:lv_res
					});
	endrule:rl_wallace_tree_part2

	rule rl_rb_nb1;
		//$display("Executing FMUL stage 2-3");
		// The Redundant Binary product generated in the previous stage is converted into the normal binary form.
		//let normal_binary_product=rb_nb(stage3.first().stage3);
		let data_from_stage3= ff_stage3.first();
		let normal_binary_product1=rb_nb1(data_from_stage3.stage3);
		//final_result<= tagged Valid (Stage4_data{final_result:normal_binary_product});
		ff_stage3.deq();
		ff_stage3a.enq(Stage3a_data{
									fsr:data_from_stage3.fsr,
				                    rounding_mode : data_from_stage3.rounding_mode,
									summed_exponent:data_from_stage3.summed_exponent,
									sign :data_from_stage3.sign,
									infinity:data_from_stage3.infinity,
									invalid:data_from_stage3.invalid,
									zero:data_from_stage3.zero,
									stage3a:{data_from_stage3.stage3,normal_binary_product1}
					});
		endrule:rl_rb_nb1
	
	rule rl_rb_nb2;
		// The Redundant Binary product generated in the previous stage is converted into the normal binary form.
		//let normal_binary_product=rb_nb(stage3.first().stage3);
		//$display("Executing FMUL stage 2-4");
		let data_from_stage3a= ff_stage3a.first();
		let data1 = data_from_stage3a.stage3a[144:17];
		let data2 = data_from_stage3a.stage3a[16:0];
		let normal_binary_product2=rb_nb2(data1,data2);
		ff_stage3b.enq (Stage3b_data{
									fsr:data_from_stage3a.fsr,
				                    rounding_mode:data_from_stage3a.rounding_mode,
									summed_exponent:data_from_stage3a.summed_exponent,
									sign :data_from_stage3a.sign,
									infinity:data_from_stage3a.infinity,
									invalid:data_from_stage3a.invalid,
									zero:data_from_stage3a.zero,
									stage3b:{data1,normal_binary_product2}
					});
		ff_stage3a.deq();
	endrule:rl_rb_nb2
	
	rule rl_rb_nb3;
		// The Redundant Binary product generated in the previous stage is converted into the normal binary form.
		//let normal_binary_product=rb_nb(stage3.first().stage3);
		let data_from_stage3b= ff_stage3b.first();
		let data1 = data_from_stage3b.stage3b[160:33];
		let data2 = data_from_stage3b.stage3b[32:0];
		let normal_binary_product3=rb_nb3(data1,data2);
		ff_stage3c.enq (Stage3c_data{
									fsr:data_from_stage3b.fsr,
				                    rounding_mode:data_from_stage3b.rounding_mode,
									summed_exponent:data_from_stage3b.summed_exponent,
									sign :data_from_stage3b.sign,
									infinity:data_from_stage3b.infinity,
									invalid:data_from_stage3b.invalid,
									zero:data_from_stage3b.zero,
									stage3c:{data1,normal_binary_product3}
					});
		ff_stage3b.deq();
		//$display("Executing FMUL stage 2-5. Data=%h",normal_binary_product3);
	endrule:rl_rb_nb3
	
	rule rl_rb_nb4;
		// The Redundant Binary product generated in the previous stage is converted into the normal binary form.
		//let normal_binary_product=rb_nb(stage3.first().stage3);
		let lv_data_from_stage3c= ff_stage3c.first();
		let data1 = lv_data_from_stage3c.stage3c[176:49];
		let data2 = lv_data_from_stage3c.stage3c[48:0];
		let normal_binary_product4=rb_nb4(data1,data2);
		ff_final_result.enq(Stage4_data{
									fsr:lv_data_from_stage3c.fsr,
				                    rounding_mode:lv_data_from_stage3c.rounding_mode,
									summed_exponent:lv_data_from_stage3c.summed_exponent,
									sign : lv_data_from_stage3c.sign,
									infinity:lv_data_from_stage3c.infinity,
									zero:lv_data_from_stage3c.zero,
									invalid:lv_data_from_stage3c.invalid,
									final_result:normal_binary_product4
						});
		//$display("Executing FMUL stage 2-6. Output=%h",normal_binary_product4);
		ff_stage3c.deq();
	endrule:rl_rb_nb4
	//Cycle 1
	method Action _start( Bit#(32) _operand1, Bit#(32) _operand2, Bit#(32) _fsr, Bit#(3) _rounding_mode, bit _sign, Bit#(10) _summed_exponent, bit _invalid, Bit#(1) _infinity, Bit#(1) _zero);
		//$display("Executing FMUL stage 2");
		Bit#(33) lv_mult={_operand1,0};		// lv_mult		= multiplier appended with a zero, a requirement of booth's second order algorithm
		Bit#(64) lv_multp={32'b0,_operand2};	// lv_multp	= multiplicand
		// Sign Extension of the multiplicand as required by the booth's algorithm.
		if(_operand2[31]==1)
			lv_multp[63:32]='d-1;
		Bit#(64) lv_lmultp = lv_multp<<1;	// lv_lmultp	= multiplicand left shifted one bit position
			
		// Generation of the 16 partial products using Booth's second order algorithm. The i+1 i i-1 th bits are used as the select bits
		// These 16 partial products are converted into redundant binary partial products by taking two at a time.i.e every adjacent partial product.
		// To form a RB number, the two's complement of the second number is needed. So, every odd numbered partial product is inverted. To avoid an addition of 1
		// which will involve a a carry propagation, we take these 8 1's along with a 64'b0 to form the 9th partial product.
		// The last two bit positions is due to the left shifting of two bits for adjacent partial products. Since, the odd numbered partial products
		// are inverted, we append one's. For even numbered partial products, we append zeroes.
		
		Vector#(16,Bit#(64)) lv_pp = replicate(0);
		lv_pp[0][63:0]=gen_pp(lv_multp,lv_lmultp,lv_mult[2:0],0)[63:0];
		lv_pp[1][63:0]={gen_pp(lv_multp,lv_lmultp,lv_mult[4:2],1)[61:0],2'b11};
		lv_pp[2][63:2]={gen_pp(lv_multp,lv_lmultp,lv_mult[6:4],0)[59:0],2'b00};
		lv_pp[3][63:4]={gen_pp(lv_multp,lv_lmultp,lv_mult[8:6],1)[57:0],2'b11};
		lv_pp[4][63:6]={gen_pp(lv_multp,lv_lmultp,lv_mult[10:8],0)[55:0],2'b00};
		lv_pp[5][63:8]={gen_pp(lv_multp,lv_lmultp,lv_mult[12:10],1)[53:0],2'b11};
		lv_pp[6][63:10]={gen_pp(lv_multp,lv_lmultp,lv_mult[14:12],0)[51:0],2'b00};
		lv_pp[7][63:12]={gen_pp(lv_multp,lv_lmultp,lv_mult[16:14],1)[49:0],2'b11};
		lv_pp[8][63:14]={gen_pp(lv_multp,lv_lmultp,lv_mult[18:16],0)[47:0],2'b00};
		lv_pp[9][63:16]={gen_pp(lv_multp,lv_lmultp,lv_mult[20:18],1)[45:0],2'b11};
		lv_pp[10][63:18]={gen_pp(lv_multp,lv_lmultp,lv_mult[22:20],0)[43:0],2'b00};
		lv_pp[11][63:20]={gen_pp(lv_multp,lv_lmultp,lv_mult[24:22],1)[41:0],2'b11};
		lv_pp[12][63:22]={gen_pp(lv_multp,lv_lmultp,lv_mult[26:24],0)[39:0],2'b00};
		lv_pp[13][63:24]={gen_pp(lv_multp,lv_lmultp,lv_mult[28:26],1)[37:0],2'b11};
		lv_pp[14][63:26]={gen_pp(lv_multp,lv_lmultp,lv_mult[30:28],0)[35:0],2'b00};
		lv_pp[15][63:28]={gen_pp(lv_multp,lv_lmultp,lv_mult[32:30],1)[33:0],2'b11};
		
		// The 16 partial products are stored in the stage1 FIFO
		ff_stage1.enq(Stage1_data{	fsr:_fsr,
				                    rounding_mode:_rounding_mode,
									summed_exponent:_summed_exponent,
									sign :_sign,
									zero:_zero,
									infinity:_infinity,
									invalid:_invalid,
									stage1:lv_pp});
	endmethod

	method Stage4_data result_();
		return ff_final_result.first();
	endmethod

	method Action _deque();
		ff_final_result.deq();
	endmethod

endmodule:mkinteger_multiplier_for_spfmul

		/*		Test Bench 		*/
/*
(*synthesize*)
module mkTb_integer_multiplier_for_spfmul(Empty);

	Reg#(Bit#(32)) rg_clock <-mkReg(0);
	Ifc_integer_multiplier_for_spfmul be <- mkinteger_multiplier_for_spfmul();

	rule rl_increment;
		rg_clock<=rg_clock+1;
		$display("CLOCK=%d",rg_clock);

		if(rg_clock=='d20)
		$finish(0);
	endrule:rl_increment
   
	rule rl_give_input(rg_clock=='d1);
		be._start(32'd14, 32'd45, 5'd10,32'd124,32'd6500,4'd12,0,0,0,0,0);
	endrule:rl_give_input
endmodule:mkTb_integer_multiplier_for_spfmul */
endpackage:integermultiplier_for_spfpu
