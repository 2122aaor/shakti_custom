// Copyright (c) 2007--2009 Bluespec, Inc.  All rights reserved.
// $Revision: 32843 $
// $Date: 2013-12-16 16:25:57 +0000 (Mon, 16 Dec 2013) $

package AHB;

////////////////////////////////////////////////////////////////////////////////
///
////////////////////////////////////////////////////////////////////////////////

import AHBArbiter::*;
import AHBBus::*;
import AHBDefines::*;
import AHBMaster::*;
import AHBPC::*;
import AHBSlave::*;

////////////////////////////////////////////////////////////////////////////////
///
////////////////////////////////////////////////////////////////////////////////

export AHBArbiter::*;
export AHBBus::*;
export AHBDefines::*;
export AHBMaster::*;
export AHBPC::*;
export AHBSlave::*;

endpackage
