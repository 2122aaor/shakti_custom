// Copyright (c) 2007--2009 Bluespec, Inc.  All rights reserved.
// $Revision: 32843 $
// $Date: 2013-12-16 16:25:57 +0000 (Mon, 16 Dec 2013) $

package TLM;

////////////////////////////////////////////////////////////////////////////////
///
////////////////////////////////////////////////////////////////////////////////

import TLMCBusAdapter::*;
import TLMDefines::*;
import TLMRam::*;
import TLMReadWriteRam::*;
import TLMReduce::*;
import TLMUtils::*;

////////////////////////////////////////////////////////////////////////////////
///
////////////////////////////////////////////////////////////////////////////////

export TLMCBusAdapter::*;
export TLMDefines::*;
export TLMRam::*;
export TLMReadWriteRam::*;
export TLMReduce::*;
export TLMUtils::*;

endpackage
