package functions;

// this function is used to count the number of trailing zeros.
// i.e is the number of zeros before the first 1, starting from the MSB
//*************************Double precision**********************
function Bit#(11) fn_count_zeros_on_right(Bit#(57) mantissa);
	if(mantissa[0]==1)
		return 0;
	else if(mantissa[1]==1)
		return 'd1;
	else if(mantissa[2]==1)
		return 'd2;
	else if(mantissa[3]==1)
		return 'd3;
	else if(mantissa[4]==1)
		return 'd4;
	else if(mantissa[5]==1)
		return 'd5;
	else if(mantissa[6]==1)
		return 'd6;
	else if(mantissa[7]==1)
		return 'd7;
	else if(mantissa[8]==1)
		return 'd8;
	else if(mantissa[9]==1)
		return 'd9;
	else if(mantissa[10]==1)
		return 'd10;
	else if(mantissa[11]==1)
		return 'd11;
	else if(mantissa[12]==1)
		return 'd12;
	else if(mantissa[13]==1)
		return 'd13;
	else if(mantissa[14]==1)
		return 'd14;
	else if(mantissa[15]==1)
		return 'd15;
	else if(mantissa[16]==1)
		return 'd16;
	else if(mantissa[17]==1)
		return 'd17;
	else if(mantissa[18]==1)
		return 'd18;
	else if(mantissa[19]==1)
		return 'd19;
	else if(mantissa[20]==1)
		return 'd20;
	else if(mantissa[21]==1)
		return 'd21;
	else if(mantissa[22]==1)
		return 'd22;
	else if(mantissa[23]==1)
		return 'd23;
	else if(mantissa[24]==1)
		return 'd24;
	else if(mantissa[25]==1)
		return 'd25;
	else if(mantissa[26]==1)
		return 'd26;
	else if(mantissa[27]==1)
		return 'd27;
	else if(mantissa[28]==1)
		return 'd28;
	else if(mantissa[29]==1)
		return 'd29;
	else if(mantissa[30]==1)
		return 30;
	else if(mantissa[31]==1)
		return 'd31;
	else if(mantissa[32]==1)
		return 'd32;
	else if(mantissa[33]==1)
		return 'd33;
	else if(mantissa[34]==1)
		return 'd34;
	else if(mantissa[35]==1)
		return 'd35;
	else if(mantissa[36]==1)
		return 'd36;
	else if(mantissa[37]==1)
		return 'd37;
	else if(mantissa[38]==1)
		return 'd38;
	else if(mantissa[39]==1)
		return 'd39;
	else if(mantissa[40]==1)
		return 40;
	else if(mantissa[41]==1)
		return 'd41;
	else if(mantissa[42]==1)
		return 'd42;
	else if(mantissa[43]==1)
		return 'd43;
	else if(mantissa[44]==1)
		return 'd44;
	else if(mantissa[45]==1)
		return 'd45;
	else if(mantissa[46]==1)
		return 'd46;
	else if(mantissa[47]==1)
		return 'd47;
	else if(mantissa[48]==1)
		return 'd48;
	else if(mantissa[49]==1)
		return 'd49;
	else if(mantissa[50]==1)
		return 50;
	else if(mantissa[51]==1)
		return 'd51;
	else if(mantissa[52]==1)
		return 'd52;
	else if(mantissa[53]==1)
		return 'd53;
	else if(mantissa[54]==1)
		return 'd54;
	else if(mantissa[55]==1)
		return 'd55;
	else if(mantissa[56]==1)
		return 'd56;
	else return 'd0;
endfunction
//THis function is used to count the number of zeros on the left of first 1 starting from MSB 
function Bit#(6) fn_count_zeros_on_left(Bit#(56) mantissa);
	if(mantissa[55]==1)
		return 0;
	else if(mantissa[54]==1)
		return 'd1;
	else if(mantissa[53]==1)
		return 'd2;
	else if(mantissa[52]==1)
		return 'd3;
	else if(mantissa[51]==1)
		return 'd4;
	else if(mantissa[50]==1)
		return 'd5;
	else if(mantissa[49]==1)
		return 'd6;
	else if(mantissa[48]==1)
		return 'd7;
	else if(mantissa[47]==1)
		return 'd8;
	else if(mantissa[46]==1)
		return 'd9;
	else if(mantissa[45]==1)
		return 'd10;
	else if(mantissa[44]==1)
		return 'd11;
	else if(mantissa[43]==1)
		return 'd12;
	else if(mantissa[42]==1)
		return 'd13;
	else if(mantissa[41]==1)
		return 'd14;
	else if(mantissa[40]==1)
		return 'd15;
	else if(mantissa[39]==1)
		return 'd16;
	else if(mantissa[38]==1)
		return 'd17;
	else if(mantissa[37]==1)
		return 'd18;
	else if(mantissa[36]==1)
		return 'd19;
	else if(mantissa[35]==1)
		return 'd20;
	else if(mantissa[34]==1)
		return 'd21;
	else if(mantissa[33]==1)
		return 'd22;
	else if(mantissa[32]==1)
		return 'd23;
	else if(mantissa[31]==1)
		return 'd24;
	else if(mantissa[30]==1)
		return 'd25;
	else if(mantissa[29]==1)
		return 'd26;
	else if(mantissa[28]==1)
		return 'd27;
	else if(mantissa[27]==1)
		return 'd28;
	else if(mantissa[26]==1)
		return 'd29;
	else if(mantissa[25]==1)
		return 'd30;
	else if(mantissa[24]==1)
		return 'd31;
	else if(mantissa[23]==1)
		return 'd32;
	else if(mantissa[22]==1)
		return 'd33;
	else if(mantissa[21]==1)
		return 'd34;
	else if(mantissa[20]==1)
		return 'd35;
	else if(mantissa[19]==1)
		return 'd36;
	else if(mantissa[18]==1)
		return 'd37;
	else if(mantissa[17]==1)
		return 'd38;
	else if(mantissa[16]==1)
		return 'd39;
	else if(mantissa[15]==1)
		return 'd40;
	else if(mantissa[14]==1)
		return 'd41;
	else if(mantissa[13]==1)
		return 'd42;
	else if(mantissa[12]==1)
		return 'd43;
	else if(mantissa[11]==1)
		return 'd44;
	else if(mantissa[10]==1)
		return 'd45;
	else if(mantissa[9]==1)
		return 'd46;
	else if(mantissa[8]==1)
		return 'd47;
	else if(mantissa[7]==1)
		return 'd48;
	else if(mantissa[6]==1)
		return 'd49;
	else if(mantissa[5]==1)
		return 'd50;
	else if(mantissa[4]==1)
		return 'd51;
	else if(mantissa[3]==1)
		return 'd52;
	else if(mantissa[2]==1)
		return 'd53;
	else if(mantissa[1]==1)
		return 'd54;
	else if(mantissa[0]==1)
		return 'd55;
	else return 'd56;
endfunction

//*********************Single precision*********************************
function Bit#(5) fnsp_count_zeros_on_left(Bit#(27) mantissa);
	if(mantissa[26]==1)
		return 0;
	else if(mantissa[25]==1)
		return 'd1;
	else if(mantissa[24]==1)
		return 'd2;
	else if(mantissa[23]==1)
		return 'd3;
	else if(mantissa[22]==1)
		return 'd4;
	else if(mantissa[21]==1)
		return 'd5;
	else if(mantissa[20]==1)
		return 'd6;
	else if(mantissa[19]==1)
		return 'd7;
	else if(mantissa[18]==1)
		return 'd8;
	else if(mantissa[17]==1)
		return 'd9;
	else if(mantissa[16]==1)
		return 'd10;
	else if(mantissa[15]==1)
		return 'd11;
	else if(mantissa[14]==1)
		return 'd12;
	else if(mantissa[13]==1)
		return 'd13;
	else if(mantissa[12]==1)
		return 'd14;
	else if(mantissa[11]==1)
		return 'd15;
	else if(mantissa[10]==1)
		return 'd16;
	else if(mantissa[9]==1)
		return 'd17;
	else if(mantissa[8]==1)
		return 'd18;
	else if(mantissa[7]==1)
		return 'd19;
	else if(mantissa[6]==1)
		return 'd20;
	else if(mantissa[5]==1)
		return 'd21;
	else if(mantissa[4]==1)
		return 'd22;
	else if(mantissa[3]==1)
		return 'd23;
	else if(mantissa[2]==1)
		return 'd24;
	else if(mantissa[1]==1)
		return 'd25;
	else if(mantissa[0]==1)
		return 'd26;
	else return 'd0;
endfunction

function Bit#(8) fnsp_count_zeros_on_right(Bit#(28) mantissa);
	if(mantissa[0]==1)
		return 0;
	else if(mantissa[1]==1)
		return 'd1;
	else if(mantissa[2]==1)
		return 'd2;
	else if(mantissa[3]==1)
		return 'd3;
	else if(mantissa[4]==1)
		return 'd4;
	else if(mantissa[5]==1)
		return 'd5;
	else if(mantissa[6]==1)
		return 'd6;
	else if(mantissa[7]==1)
		return 'd7;
	else if(mantissa[8]==1)
		return 'd8;
	else if(mantissa[9]==1)
		return 'd9;
	else if(mantissa[10]==1)
		return 'd10;
	else if(mantissa[11]==1)
		return 'd11;
	else if(mantissa[12]==1)
		return 'd12;
	else if(mantissa[13]==1)
		return 'd13;
	else if(mantissa[14]==1)
		return 'd14;
	else if(mantissa[15]==1)
		return 'd15;
	else if(mantissa[16]==1)
		return 'd16;
	else if(mantissa[17]==1)
		return 'd17;
	else if(mantissa[18]==1)
		return 'd18;
	else if(mantissa[19]==1)
		return 'd19;
	else if(mantissa[20]==1)
		return 'd20;
	else if(mantissa[21]==1)
		return 'd21;
	else if(mantissa[22]==1)
		return 'd22;
	else if(mantissa[23]==1)
		return 'd23;
	else if(mantissa[24]==1)
		return 'd24;
	else if(mantissa[25]==1)
		return 'd25;
	else if(mantissa[26]==1)
		return 'd26;
	else if(mantissa[27]==1)
		return 'd27;
	else return 'd0;
endfunction

function Bit#(9) fn_count_leadingzeros(Bit#(56) mantissa);
	if(mantissa[55]==1)
		return 0;
	else if(mantissa[54]==1)
		return 1;
	else if(mantissa[53]==1)
		return 2;
	else if(mantissa[52]==1)
		return 3;
	else if(mantissa[51]==1)
		return 4;
	else if(mantissa[50]==1)
		return 5;
	else if(mantissa[49]==1)
		return 6;
	else if(mantissa[48]==1)
		return 7;
	else if(mantissa[47]==1)
		return 8;
	else if(mantissa[46]==1)
		return 9;
	else if(mantissa[45]==1)
		return 10;
	else if(mantissa[44]==1)
		return 11;
	else if(mantissa[43]==1)
		return 12;
	else if(mantissa[42]==1)
		return 13;
	else if(mantissa[41]==1)
		return 14;
	else if(mantissa[40]==1)
		return 15;
	else if(mantissa[39]==1)
		return 16;
	else if(mantissa[38]==1)
		return 17;
	else if(mantissa[37]==1)
		return 18;
	else if(mantissa[36]==1)
		return 19;
	else if(mantissa[35]==1)
		return 20;
	else if(mantissa[34]==1)
		return 21;
	else if(mantissa[33]==1)
		return 22;
	else if(mantissa[32]==1)
		return 23;
	else if(mantissa[31]==1)
		return 24;
	else if(mantissa[30]==1)
		return 25;
	else if(mantissa[29]==1)
		return 26;
	else if(mantissa[28]==1)
		return 27;
	else if(mantissa[27]==1)
		return 28;
	else if(mantissa[26]==1)
		return 29;
	else if(mantissa[25]==1)
		return 30;
	else if(mantissa[24]==1)
		return 31;
	else if(mantissa[23]==1)
		return 32;
	else if(mantissa[22]==1)
		return 33;
	else if(mantissa[21]==1)
		return 34;
	else if(mantissa[20]==1)
		return 35;
	else if(mantissa[19]==1)
		return 36;
	else if(mantissa[18]==1)
		return 37;
	else if(mantissa[17]==1)
		return 38;
	else if(mantissa[16]==1)
		return 39;
	else if(mantissa[15]==1)
		return 40;
	else if(mantissa[14]==1)
		return 41;
	else if(mantissa[13]==1)
		return 42;
	else if(mantissa[12]==1)
		return 43;
	else if(mantissa[11]==1)
		return 44;
	else if(mantissa[10]==1)
		return 45;
	else if(mantissa[9]==1)
		return 46;
	else if(mantissa[8]==1)
		return 47;
	else if(mantissa[7]==1)
		return 48;
	else if(mantissa[6]==1)
		return 49;
	else if(mantissa[5]==1)
		return 50;
	else if(mantissa[4]==1)
		return 51;
	else if(mantissa[3]==1)
		return 52;
	else if(mantissa[2]==1)
		return 53;
	else if(mantissa[1]==1)
		return 54;
	else if(mantissa[0]==1)
		return 55;
	else 
		return 0;
	
endfunction
	
endpackage
