// Copyright (c) 2007--2009 Bluespec, Inc.  All rights reserved.
// $Revision: 32843 $
// $Date: 2013-12-16 16:25:57 +0000 (Mon, 16 Dec 2013) $

package Axi;

////////////////////////////////////////////////////////////////////////////////
///
////////////////////////////////////////////////////////////////////////////////

import AxiDefines::*;
import AxiMaster::*;
import AxiSlave::*;
import AxiRdBus::*;
import AxiWrBus::*;
import AxiPC::*;
import AxiMonitor::*;

////////////////////////////////////////////////////////////////////////////////
///
////////////////////////////////////////////////////////////////////////////////

export AxiDefines::*;
export AxiMaster::*;
export AxiSlave::*;
export AxiRdBus::*;
export AxiWrBus::*;
export AxiPC::*;
export AxiMonitor::*;

endpackage
