`define REG_WIDTH 64
`define PRF_SIZE 128
