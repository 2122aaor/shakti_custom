// Copyright (c) 2007--2009 Bluespec, Inc.  All rights reserved.
// $Revision: 32843 $
// $Date: 2013-12-16 16:25:57 +0000 (Mon, 16 Dec 2013) $

package TLM2;

////////////////////////////////////////////////////////////////////////////////
///
////////////////////////////////////////////////////////////////////////////////

import TLM2BRAM::*;
import TLM2CBusAdapter::*;
import TLM2Defines::*;
import TLM2Ram::*;
import TLM2ReadWriteRam::*;
import TLM2Reduce::*;
import TLM2Utils::*;
import BusSwitch::*;

////////////////////////////////////////////////////////////////////////////////
///
////////////////////////////////////////////////////////////////////////////////

export TLM2BRAM::*;
export TLM2CBusAdapter::*;
export TLM2Defines::*;
export TLM2Ram::*;
export TLM2ReadWriteRam::*;
export TLM2Reduce::*;
export TLM2Utils::*;
export BusSwitch::*;

endpackage
